`include "../define.v"

module exu (

);
    
endmodule