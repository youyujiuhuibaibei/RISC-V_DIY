`include "../define.v"

module cpu_top (
    input clk,
    input rst_n
);




endmodule