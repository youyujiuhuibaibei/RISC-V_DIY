`include "../define.v"
//`include "cpu_top.v"
`include "Data_mem.v"
`include "Inst_mem.v"
`include "ifu.v"
`include "if_id.v"
`include "idu.v"
`include "id_ex.v"
`include "exu.v"
`include "ex_mem.v"
`include "memu.v"
`include "mem_wb.v"
`include "wbu.v"
`include "regs.v"