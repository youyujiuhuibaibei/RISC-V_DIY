`include "../define.v"

module cpu_top (
    input clk,
    input rst_n
);

wire [31:0] PC;
wire [31:0] Inst_in;
wire [31:0] Inst_out;




endmodule